library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package MyDef is
    constant n:integer:=16;
end package MyDef;